-- Fichero MEDTH.vhd
-- Modelo VHDL 2002 del nivel superior de la jerarquia del circuito medidor de temperatura y humedad relativa

-- Especificacion: MEMTEMP posee interfaces con un teclado hexadecimal, un sensor de temperatura y humedad y 8 displays
-- de 7 segmentos. Ademas, posee un reloj que indica horas, minutos y segundos. El sistema realiza lecturas de humedad
-- relativa y temperatura cada 0.5 seg. Mediante el teclado hexadecimal es posible configurar la presentacion de esta
-- informacion en 4 modos: solo reloj, solo temperatura, solo humedad y todo; en este ultimo modo la informacion se
-- presenta secuencialmente (reloj, temperatura, humedad, reloj...) y cada dato se introduce por la izquierda de la
-- barra de displays de manera semejante a la que se utiliza en los visualizadores comerciales (p. ej, en farmacias).
-- El reloj tiene dos modos de funcionamiento (12 y 24 hs) y la hora puede programarse, todo ello utilizando tambien
-- el teclado hexadecimal.

-- Este modelo es estructural y contiene los siguientes bloques funcionales:

-- 1.- CTRL_TEC:    Controlador de teclado hexadecimal. Genera la tecla pulsada y una segnal de habilitacion
--                  cada vez que se pulsa una de las teclas del teclado.
-- 2.- RELOJ_12_24: Reloj con formato 12-24. Reloj programable que muestra horas, minutos y segundos. La programacion
--                  puede realizarse con el teclado hexadecimal.
-- 3.- TIMER:       Temporizador que genera tics de 5 ms, 250ms y 1s, necesaros para el funcionamiento de los
--                  otros modulos.
-- 4.- I2C:         Controlador I2C. Interfaz I2C bidireccional.
-- 5.- DISPLAY:     Controlador de displays de 7 segmentos. Gestiona la presentacion de la temperatura, humedad relativa 
--                  y el reloj. Posee 4 modos de trabajo que pueden configurarse con el teclado hexadecimal.
-- 6.- THPROC:      Procesador de temperatura y humedad. Maneja al controlador I2C para que realice lecturas
--                  periodicas de temperatura y humedad relativa y genera valores BCD listos para ser presentados
--                  en los displays.
-- 7.- PLL:         PLL que genera el reloj de 100 MHz a partir del reloj de 50 MHz de la tarjeta DECA-MAX10
--
--    Designer: DTE
--    Version: 1.0
--    Fecha: 01-01-2017


library ieee;
use ieee.std_logic_1164.all;

entity MEDTH is 
generic(                        -- Los valores por defecto para sintesis logica. En la simulacion se utilizan otros valores para escalarla
    DIV_125ms : natural := 24;
    DIV_1ms : natural := 99999;
    TICS_2s : natural := 400;
    PLL_ARCH: string :="syn"
   );
port(
    clk           : in std_logic;
    nRst          : in std_logic;
    SDA           : inout  std_logic;
    SCL           : inout  std_logic
    );  
end entity;

architecture struct of MEDTH is
  signal clk_100:        std_logic;
  signal tic_1ms:        std_logic;
  signal tic_5ms:        std_logic;
  signal tic_125ms:      std_logic;
  signal tic_025s:       std_logic;
  signal tic_1s:         std_logic;
  signal rd:             std_logic;
  signal we:             std_logic;
  signal add:            std_logic_vector(1 downto 0);
  signal dato_in:        std_logic_vector(7 downto 0);  
  signal dato_out:       std_logic_vector(7 downto 0);
  
begin

TIMER: entity work.timer(rtl) 
generic map(
    DIV_125ms   => DIV_125ms,
    DIV_1ms     => DIV_1ms
    )
port map(
    clk         => clk_100,
    nRst        => nRst,
    tic_125ms   => tic_125ms,
    tic_025s    => tic_025s,
    tic_1s      => tic_1s,
    tic_5ms     => tic_5ms,
    tic_1ms     => tic_1ms
    );
I2C: entity work.periferico_i2c(estructural) port map(
     clk        => clk_100,
     nRst       => nRst,
     we         => we,
     rd         => rd,
     add        => add,
     dato_in    => dato_in,
     dato_out   => dato_out,               
     SDA        => SDA,                    
     SCL        => SCL                    
    );
	
THPROC: entity work.procesador_medida(rtl) port map(
     clk         => clk_100,
     nRst        => nRst,
     tic_0_25s   => tic_025s,
     we          => we,
     rd          => rd,
     add         => add,
     dato_w      => dato_in,
     dato_r      => dato_out,
     dato_leido  => open
    );

sintesis: if PLL_ARCH = "syn" generate
PLL: entity work.pll_100mhz(syn) port map( 
     inclk0      => clk,
     c0          => clk_100
    );	
end generate sintesis;

simulacion: if PLL_ARCH = "sim" generate
PLL: entity work.pll_100mhz(sim) port map( 
     inclk0      => clk,
     c0          => clk_100
    );	
end generate simulacion;
assert(PLL_ARCH="syn" or PLL_ARCH="sim")
report"No se ha definido ninguna arquitectura para el PLL"
severity failure;
end struct;